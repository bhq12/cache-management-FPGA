----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:10:36 10/05/2016 
-- Design Name: 
-- Module Name:    cache_controller_frog - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cache_controller_frog is
	port(data_in, data_from_device, address_in: in std_logic_vector(7 downto 0);
	operation : in std_logic_vector(1 downto 0);
	data_to_device : out std_logic_vector(7 downto 0);
	data_result : out std_logic_vector(7 downto 0);
	address_out : out std_logic_vector(7 downto 0);
	rw_out : out std_ulogic;
	hm : in std_ulogic; --hit/miss
	em, ec : out std_ulogic; -- enable main/cache
	read_ready : in std_ulogic);
end cache_controller_frog;

architecture Behavioral of cache_controller_frog is

begin
	process
	begin
		if operation = "00" then
			address_out <= address_in;
			data_to_device <= data_in;
			data_result <= data_from_device;
			ec <= '1';
		end if;
		
--		if operation = "11" then
--
--		end
		
		if operation = "01" then
			rw_out <= '1'; -- read
		end if;
		
		if operation = "01" then
			rw_out <= '0'; -- write
		end if;
		
		if rising_edge(hm) then
			--miss has occurred
			em <= '1';--enable main memory
			ec <= '0';--disable cache
		end if;
		
		if rising_edge(read_ready) then
			data_to_device <= data_from_device;
			rw_out <= '0'; --write
			ec <= '1';
			em <= '0';
		end if;
	end process;
end Behavioral;